///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File Name: apb_mstr_driver.sv
// Description: APB Master driver
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class apb_master_driver extends uvm_driver#(apb_seq_item);
    `uvm_component_utils(apb_master_driver)
    
  
  
  
  // virtual interface instance
  virtual apb_interface   apb_intf_drv;
  
  
  // analysis port declaration
  uvm_analysis_port#(apb_seq_item) drv2scb;
    
    
    
    // constructor function
  function new(string name="apb_master_driver", uvm_component parent=null);
    super.new(name, parent);
    // create the analysis port
    drv2scb = new("drv2scb", this);
        
  endfunction: new
    
    // build_phase
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    
    if(!uvm_config_db#(virtual apb_interface)::get(this, "", "apb_interface", apb_intf_drv)) begin
      `uvm_fatal("NO APB_INTF ERROR", "driver cannot obtain virtual interface! please check config_db setting")
    end
    
  endfunction: build_phase
    
    // connect_phase
  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
  endfunction: connect_phase
    
    // run_phase
  virtual task run_phase(uvm_phase phase);
  	apb_seq_item item;
        
  // reset the interface
    apb_intf_drv.reset_intf();
        
        // get data from sequencer and drive to DUT
        forever begin
          @(apb_intf_drv.cb);
          seq_item_port.get_next_item(item);
          if(item.op_type == WRITE) begin
            wr_data(item);
            // write expected data to analysis port
            drv2scb.write(item);
          end
          else if(item.op_type == READ) begin
            rd_data(item);
          end
          seq_item_port.item_done();
        end    
  endtask: run_phase
  /*
    Inheritance
    uvm_driver (Base class): Has already declared and instantiated seq_item_port.
    my_driver (Derived class): Directly uses seq_item_port, no need to redeclare.
 */
    
    ////////////////////////////////////////////////////////////////////
    // task name: wr_data
    // input parameter: apb_seq_item
    // Description: write data to dut
    ////////////////////////////////////////////////////////////////////
  task wr_data(input apb_seq_item item);
        apb_intf_drv.cb.PSEL <= 1;
        apb_intf_drv.cb.PWRITE <= 1;
        apb_intf_drv.cb.PADDR <= item.ADDR;
        apb_intf_drv.cb.PWDATA <= item.DATA;
        apb_intf_drv.cb.PENABLE <= 0;
        @(apb_intf_drv.cb);
        apb_intf_drv.cb.PENABLE <= 1;
        @(apb_intf_drv.cb);
        wait(apb_intf_drv.cb.PREADY == 1);
        apb_intf_drv.cb.PENABLE <= 0;
        apb_intf_drv.cb.PSEL <= 0;
        @(apb_intf_drv.cb);
  endtask: wr_data
    
    ////////////////////////////////////////////////////////////////////
    // task name: rd_data
    // input parameter: addr, data
    // Description: read data to dut 
	// I modify github code by add a damn clk for data of odd address 
    ////////////////////////////////////////////////////////////////////
  task rd_data(input apb_seq_item item);
        apb_intf_drv.cb.PSEL <= 1;
        apb_intf_drv.cb.PWRITE <= 0;
        apb_intf_drv.cb.PADDR <= item.ADDR;
        apb_intf_drv.cb.PENABLE <= 0;
        @(apb_intf_drv.cb);
        apb_intf_drv.cb.PENABLE <= 1;
    	@(apb_intf_drv.cb);
        wait(apb_intf_drv.cb.PREADY == 1);
        apb_intf_drv.cb.PENABLE <= 0;
        apb_intf_drv.cb.PSEL <= 0;
    	@(apb_intf_drv.cb);
  endtask: rd_data
endclass: apb_master_driver